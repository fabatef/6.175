import ProcTypes::*;
import MemTypes::*;
import Types::*;
import CacheTypes::*;
import MessageFifo::*;
import Vector::*;
import FShow::*;

// TODO: implement parent protocol processor

module mkPPP(MessageGet c2m, MessagePut m2c, WideMem mem, Empty ifc);

endmodule

