import CacheTypes::*;
import Vector::*;
import MemTypes::*;
import Types::*;
import ProcTypes::*;
import Fifo::*;
import Ehr::*;

// TODO
module mkICache(WideMem mem, ICache ifc);

endmodule

